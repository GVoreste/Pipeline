package Pipeline is
    


end Pipeline;

package body Pipeline is
end Pipeline;